* EESchema Netlist Version 1.1 (Spice format) creation date: Tue 04 Aug 2015 19:43:35 BST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

*Sheet Name:/
R1  +5V N-000003 10K		
SW1  GND N-000003 REED		
R2  N-000003 ? 10K		

.end
